module rule_ram 
#(parameter DATA_WIDTH = 32
)
(
	input [4:0] addr_r,
	input [4:0] addr_w,
	input [DATA_WIDTH-1:0] din,
	output [DATA_WIDTH-1:0] dout,
	input we,
	input clk
);




endmodule 
